----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:50:55 12/30/2016 
-- Design Name: 
-- Module Name:    inst_motor_ascensor - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity inst_motor_ascensor is
    Port ( accionar_ascensor : in  STD_LOGIC;
           actuador_motor_subir : out  STD_LOGIC;
           actuador_motor_bajar : out  STD_LOGIC);
end inst_motor_ascensor;

architecture Behavioral of inst_motor_ascensor is

begin


end Behavioral;

